module noise_gen ();

endmodule