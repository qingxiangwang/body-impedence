module dpsd_simu(dds_noise_filter_out,clk);

 output dds_noise_filter_out;
 input clk;
 input noise;

always @(posedge clk) begin
  a =0;
  end
endmodule