module dds (sin_wave,system_clk,FT_Word);



output sin_wave;
input system_clk;
input FT_Word;
endmodule

//---------------------------------------------
//


