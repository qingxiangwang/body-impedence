module dpsd_simu(output reg a,input clk);
always @(posedge clk) begin
  a =0;
  end
endmodule